`timescale 1ns / 1ps

module npu_top_tb;

    reg clk = 0;
    reg rst = 1;
    reg [63:0] image;
    wire [15:0] logit0, logit1, logit2, logit3, logit4;
    wire [15:0] logit5, logit6, logit7, logit8, logit9;
    wire done;
    wire [3:0] predict_idx;

    npu_top dut (
        .clk(clk),
        .rst(rst),
        .image(image),
        .logit0(logit0), .logit1(logit1), .logit2(logit2), .logit3(logit3), .logit4(logit4),
        .logit5(logit5), .logit6(logit6), .logit7(logit7), .logit8(logit8), .logit9(logit9),
        .done(done), .predict_idx(predict_idx)
    );

    always #10 clk = ~clk;

    // === Memory holding 256 test images ===
    reg [63:0] image_mem [0:255];      // 256 images, each 64-bit
    reg [3:0]  predict_result [0:255]; // store predicted class index

    initial begin
        image_mem[0] = 64'b0001110000110000001000000010000000111100001101000011110000001100;  // Label: 9
image_mem[1] = 64'b0001110000100100001000000011000000011000000100000001010000011000;  // Label: 3
image_mem[2] = 64'b0000100000011000000100000001000000100100010001000111110001111000;  // Label: 7
image_mem[3] = 64'b0011110001100100000001000000110000011000000100000001110000011100;  // Label: 2
image_mem[4] = 64'b1111110000111100000110000001100000001100000011100000110000001100;  // Label: 1
image_mem[5] = 64'b0001110000011000000100000001110000001100000001100011110001111000;  // Label: 5
image_mem[6] = 64'b0110100000111000000100000001000000100000001001000010110000011000;  // Label: 2
image_mem[7] = 64'b0000110000011000000100000001110000001100000001000000110000111100;  // Label: 5
image_mem[8] = 64'b0000110000111100001110000001000000010000000100000001110000001100;  // Label: 2
image_mem[9] = 64'b0011100000011000000110000001100000010000000110000011100000011000;  // Label: 1
image_mem[10] = 64'b0011000000100000001000000011110000110100011001000110100001100000;  // Label: 9
image_mem[11] = 64'b0000100000001000000111000111111000110100000101000000110000001000;  // Label: 4
image_mem[12] = 64'b0001100000111100001001000000000000000000001001000011110000011000;  // Label: 0
image_mem[13] = 64'b0001100000010000001111000111011001100100010011000000100000010000;  // Label: 4
image_mem[14] = 64'b0000110000111100000111000001000000010000001100000001110000011100;  // Label: 2
image_mem[15] = 64'b0011110000101000001000000011100000011000000100000011110000011000;  // Label: 3
image_mem[16] = 64'b0000100000011000000100000011110000110000001000000110100001111000;  // Label: 7
image_mem[17] = 64'b0011100000101000001010000011100000011100001001000010110000111000;  // Label: 8
image_mem[18] = 64'b0001110000100100001011000001100000111100000101000000110000001100;  // Label: 8
image_mem[19] = 64'b0001000000010000001111000011110000010100001010000001100000010000;  // Label: 4
image_mem[20] = 64'b0001110000110000001100000001000000010000001100000011110000111100;  // Label: 3
image_mem[21] = 64'b0001110000110000001100000011000000111100001111100011110000001100;  // Label: 9
image_mem[22] = 64'b0000010000001000000011000011110000110000001000000011100000111000;  // Label: 7
image_mem[23] = 64'b0001100000011000000100000001100000001110000011100000110000111000;  // Label: 5
image_mem[24] = 64'b0011100001101100001111000000010000000100000001000000110000001000;  // Label: 6
image_mem[25] = 64'b0011100001101100011000000011000000010000000101100010110000011000;  // Label: 3
image_mem[26] = 64'b0001110000011000000110000001100000001100000011000001110000111100;  // Label: 5
image_mem[27] = 64'b0011100001100100011001000011110000000100000001000000110000001000;  // Label: 6
image_mem[28] = 64'b0011110001100100011001000010000000111000000100000001000000011100;  // Label: 3
image_mem[29] = 64'b0001000000111110001111100010011000000100000010000001100000010000;  // Label: 4
image_mem[30] = 64'b0011100001101100011000000010000000111000001001000011110000011000;  // Label: 9
image_mem[31] = 64'b1111100000111100001000000001000000011000000110000000100000001000;  // Label: 1
image_mem[32] = 64'b0001000000011100001111100110011000000100000011000001100000011000;  // Label: 4
image_mem[33] = 64'b0001100000011000000100000011110001100100010001000000110000011000;  // Label: 4
image_mem[34] = 64'b0111100001101100001001000011110000001100000011000001110000011000;  // Label: 6
image_mem[35] = 64'b0011100000100000001000000010000000101100001101000011010000001000;  // Label: 9
image_mem[36] = 64'b0001100000010000000111000111011000110100000011000000100000010000;  // Label: 4
image_mem[37] = 64'b0000010000000100000010000001110001111000001100000011000000111100;  // Label: 7
image_mem[38] = 64'b0111000001101000011011000001110000000100000011000000100000011000;  // Label: 6
image_mem[39] = 64'b0011000001001100010011000011110000000100000011000000100000011000;  // Label: 6
image_mem[40] = 64'b0011100000110000001000000010000000111000001111000001110000001000;  // Label: 9
image_mem[41] = 64'b0011100000011100000111000001110000011100000111000001110000011000;  // Label: 1
image_mem[42] = 64'b0001110000100100001000000010000000011000000100000011010000011000;  // Label: 3
image_mem[43] = 64'b0001100000111100001111000000110000000100000011000000100000001000;  // Label: 6
image_mem[44] = 64'b0011100000111000001110000001100000111100001111000011100000110000;  // Label: 1
image_mem[45] = 64'b0001110000100000001000000011000000011000000100000001010000011100;  // Label: 3
image_mem[46] = 64'b0001110000110100001001000010010000100100001001000001110000001100;  // Label: 0
image_mem[47] = 64'b0011100001000100010011000011110000000100000001000000110000011000;  // Label: 6
image_mem[48] = 64'b0001110000100100001000000001100000001110000001000000110000111100;  // Label: 5
image_mem[49] = 64'b0001100000011000000000000011010000011100000001000111110001110000;  // Label: 5
image_mem[50] = 64'b0011100000011100001110000001110000111000000111000011100000001000;  // Label: 1
image_mem[51] = 64'b0111000001000100010000000010000000110100000100000001010000010000;  // Label: 9
image_mem[52] = 64'b0001110000011000000100000001110000001100000001000011110000111100;  // Label: 5
image_mem[53] = 64'b0011100000100000000001000011110000000100000001000001110000011000;  // Label: 6
image_mem[54] = 64'b0011100000100100000001000000010000000100000001000011110000011000;  // Label: 0
image_mem[55] = 64'b0111100001110000011000000010000000111000000111000001110000001100;  // Label: 9
image_mem[56] = 64'b0000100000011100001111000000010000000100001001000011110000001100;  // Label: 0
image_mem[57] = 64'b0011100000100100000001000000010000000100001001000010010000011000;  // Label: 0
image_mem[58] = 64'b0011000000010000000100000001000000010100000111000011100000010000;  // Label: 1
image_mem[59] = 64'b0000110000011100001100000010000000000000000001000010110000011100;  // Label: 0
image_mem[60] = 64'b0001000000010000001111000111111000110100001011000001100000010000;  // Label: 4
image_mem[61] = 64'b0001100000110000001000000010110000111100000011000000110000111000;  // Label: 5
image_mem[62] = 64'b0011100001111100000110000001000000010100000101100001110000001100;  // Label: 2
image_mem[63] = 64'b0001000000110000001111100011111000100100000011000001100000010000;  // Label: 4
image_mem[64] = 64'b0001110000100000000000000010000000011100000001000000110000111100;  // Label: 5
image_mem[65] = 64'b0000100000001000000111000011110000010010000101000010110000111000;  // Label: 7
image_mem[66] = 64'b0001100000100100001001000010010000101100001011000011110000001000;  // Label: 0
image_mem[67] = 64'b0000110000001000000110000111110000110000000100100011111000011000;  // Label: 7
image_mem[68] = 64'b0001100000100000001000000010110000111100000001000000100000111000;  // Label: 5
image_mem[69] = 64'b0001100000100000011000000111100000100100001001000011110000011000;  // Label: 9
image_mem[70] = 64'b0011110001100100010000000010000000111100000001000000010000011100;  // Label: 5
image_mem[71] = 64'b0011100000100000001000000011110000000110000001000000110000111000;  // Label: 5
image_mem[72] = 64'b0000100000001000000011000011111000110110001101000000110000001000;  // Label: 4
image_mem[73] = 64'b0000100000001000000010000111110000010000001101000011110000111000;  // Label: 7
image_mem[74] = 64'b0001100000111100001001000000010000000100001001000010110000001000;  // Label: 0
image_mem[75] = 64'b0010000000100000001111100011110001101000000100000001000000100000;  // Label: 4
image_mem[76] = 64'b0001110000011100000110000000110000001100000001000011110000011100;  // Label: 5
image_mem[77] = 64'b0001100000100100001000000000000000111100000001000000010000111000;  // Label: 5
image_mem[78] = 64'b0001110000100100000000000000000000101000001101000011010000011100;  // Label: 9
image_mem[79] = 64'b0011100000101100001000000010100000111100001101000011110000011000;  // Label: 9
image_mem[80] = 64'b0001100000110100001001000010010000100100001111000011110000001000;  // Label: 0
image_mem[81] = 64'b0000110001111100000010000001100000010000000100000000111000001100;  // Label: 2
image_mem[82] = 64'b0001110000110000001100000001000000110000001000000110010000111000;  // Label: 3
image_mem[83] = 64'b0011100001101100001001000001110000011100001001000010010000111000;  // Label: 8
image_mem[84] = 64'b0001100000110100001001000000010000100100001001000011110000011000;  // Label: 0
image_mem[85] = 64'b0111000001001000010011000010110000001100000011000000100000011000;  // Label: 6
image_mem[86] = 64'b0001100000011000001110000011111001111100000011000000100000011000;  // Label: 4
image_mem[87] = 64'b0001000000010000000111000011110001100100000001000000100000010000;  // Label: 4
image_mem[88] = 64'b0011100000110000001000000010000000110000001111000011110000011000;  // Label: 9
image_mem[89] = 64'b0001000000011000000110000001000000011110000111000011100000110000;  // Label: 1
image_mem[90] = 64'b0111100000001000000010000001000000010000000001000001110000011000;  // Label: 2
image_mem[91] = 64'b0111000000100100001011000001100000011000001010000011100000110000;  // Label: 8
image_mem[92] = 64'b0001100000111000001000000011000000011000001100000011110000111000;  // Label: 3
image_mem[93] = 64'b0011110000000100001000000010000000110100000111000000010000111100;  // Label: 5
image_mem[94] = 64'b0110100001111000000100000001000000010000000101000001110000001000;  // Label: 2
image_mem[95] = 64'b0011100000100000001000000010000000111100001000100010010000011000;  // Label: 9
image_mem[96] = 64'b0001100000111000001111000010010000100100001011000011100000011000;  // Label: 0
image_mem[97] = 64'b0001100000010000001100000011110000100100000001000000110000011000;  // Label: 4
image_mem[98] = 64'b0000100000001000000111100111111000010100001101000000110000001000;  // Label: 4
image_mem[99] = 64'b0001000000010000001111000111110000011100000110000001000000110000;  // Label: 4
image_mem[100] = 64'b0001110000100000001000000011000000011000001100000110110000111100;  // Label: 3
image_mem[101] = 64'b0000110000011000001000000010010000111100000001000000010000111000;  // Label: 5
image_mem[102] = 64'b0001100000011000001000000011000000110000001100000011110000111000;  // Label: 3
image_mem[103] = 64'b0010000000110000001100000011000000111100001110000111000000100000;  // Label: 1
image_mem[104] = 64'b0001110000110000000110000000110000011000001100000111000000111100;  // Label: 3
image_mem[105] = 64'b0000110000011000000100000001110000001110000001000000110000111100;  // Label: 5
image_mem[106] = 64'b0001000000010000000100000001110000111100011011000111100001110000;  // Label: 9
image_mem[107] = 64'b0001000000011000001111100011010000110100001110000001100000010000;  // Label: 4
image_mem[108] = 64'b1111100001111000000100000001000000110000000101100001111000011000;  // Label: 2
image_mem[109] = 64'b0001100000011000000100000011100001110000011000000111100001111000;  // Label: 7
image_mem[110] = 64'b0000100000001000000110000011110000110000001100000011100000111000;  // Label: 7
image_mem[111] = 64'b0000100000011000000111000011010000010100001001000000100000011000;  // Label: 4
image_mem[112] = 64'b0001100000011000001111100011011000010100000011000000100000011000;  // Label: 4
image_mem[113] = 64'b0011000000110000001110000001110000011100000111000011100000010000;  // Label: 1
image_mem[114] = 64'b0001110000100000001000000010000000110000001101000011010000011100;  // Label: 9
image_mem[115] = 64'b0011100000001100000011000001100000100000001010000011100000010000;  // Label: 2
image_mem[116] = 64'b0000010000001000000010000011100000010000000101000011110001101000;  // Label: 7
image_mem[117] = 64'b0001100000000100001001000001110000100100001000000010010000010000;  // Label: 8
image_mem[118] = 64'b0000100000010000000100000011110001111000011000000111100000111000;  // Label: 7
image_mem[119] = 64'b0111110000111100000010000001000000010000000100100001111000011100;  // Label: 2
image_mem[120] = 64'b0011100001101100011001000011110000000100000001000000110000011000;  // Label: 6
image_mem[121] = 64'b0001110000110000001000000010000000100100001001000000010000011100;  // Label: 9
image_mem[122] = 64'b0001000000100000001000000011111001001100010010000000100000010000;  // Label: 4
image_mem[123] = 64'b0011100001101000010001000100010000000000001000100000101000010000;  // Label: 0
image_mem[124] = 64'b0000010000001000000010000011110000010000000100000001010000011000;  // Label: 7
image_mem[125] = 64'b0011110000101100000001000000110000001000000100000001110000011100;  // Label: 2
image_mem[126] = 64'b0000100000001000001111000011100000110000001000000011110000111000;  // Label: 7
image_mem[127] = 64'b0000110000011100000110000001100000001100000001100010111000111100;  // Label: 5
image_mem[128] = 64'b0011000000101000000101000001110000011000001010000010100000110000;  // Label: 8
image_mem[129] = 64'b0000011000000100000011000011110000011000000101000011110000011100;  // Label: 7
image_mem[130] = 64'b0000110000011000001100000010000000111100000001100000010000111100;  // Label: 5
image_mem[131] = 64'b0000100000001000000110000111100000010000000101000011110000111000;  // Label: 7
image_mem[132] = 64'b0001000000010000000100000011000000100100001001000011110000110000;  // Label: 7
image_mem[133] = 64'b0001100000110100001001000010000000000100000011000011110000001000;  // Label: 0
image_mem[134] = 64'b0011100001001100011011000011110000000100000001000000110000011000;  // Label: 6
image_mem[135] = 64'b0011100001101100011011000000110000001100000011000000110000001000;  // Label: 6
image_mem[136] = 64'b0001100000010000001110000011010000100100000011000001100000010000;  // Label: 4
image_mem[137] = 64'b0111000001111100000110000001000000010000000101000001110000011000;  // Label: 2
image_mem[138] = 64'b0001100000010100000101000001110000011100001111000011110000011000;  // Label: 8
image_mem[139] = 64'b0001100000111100010001000100010000000100001011000001100000011000;  // Label: 0
image_mem[140] = 64'b0011100000100000001000000010000000111100001101000001010000011000;  // Label: 9
image_mem[141] = 64'b0001000000010000000111000111111000010100000110000001100000010000;  // Label: 4
image_mem[142] = 64'b0011100001101100010001000010010000000100000001000000110000001000;  // Label: 6
image_mem[143] = 64'b0001100000111000001000000011100000111100001001000001110000001000;  // Label: 9
image_mem[144] = 64'b0001000000110000001000000010000000111100011001000100100001110000;  // Label: 9
image_mem[145] = 64'b0001100000100100010011000011110000000100000001000000010000001000;  // Label: 6
image_mem[146] = 64'b0011100001100000010000000110000000111000001111000010010000011000;  // Label: 9
image_mem[147] = 64'b0011100000101000001001000000000000000100001001000010110000011000;  // Label: 0
image_mem[148] = 64'b0001100001110000011000000011000000011100000111000001100000011000;  // Label: 3
image_mem[149] = 64'b0001100000100000001000000011000000001110000001100000110000110000;  // Label: 5
image_mem[150] = 64'b0011100001101100001111000000110000000100000011000001110000011000;  // Label: 6
image_mem[151] = 64'b0011000000111100011011000011110000001100000011000001110000010000;  // Label: 6
image_mem[152] = 64'b0011100000100100000001000000010000100100001001000001110000011100;  // Label: 0
image_mem[153] = 64'b0011100001101100010011000011110000001100000011000000100000001000;  // Label: 6
image_mem[154] = 64'b0001100000011000000111100111011000110100001001000000100000011000;  // Label: 4
image_mem[155] = 64'b0111100001001000011000000001000000010000000101100011110000010000;  // Label: 3
image_mem[156] = 64'b0011110001100000001000000010000000111000001111000001110000001100;  // Label: 9
image_mem[157] = 64'b0011110000100000001000000011000000011000000100000011010000011100;  // Label: 3
image_mem[158] = 64'b0000100000001000000010000001100000011100001111000011110000011000;  // Label: 9
image_mem[159] = 64'b0000100000001000000111000011110000110000001100000011110000011000;  // Label: 7
image_mem[160] = 64'b0011110000100110000011000000100000011000000100000001110000001100;  // Label: 2
image_mem[161] = 64'b0011110000100100000000000010000000100000001111000011010000011100;  // Label: 9
image_mem[162] = 64'b0001100000011100001001000010010000100100001001000011110000011000;  // Label: 0
image_mem[163] = 64'b0011000000111100001101000010010001001100000010000001100000110000;  // Label: 4
image_mem[164] = 64'b0000110000010000000100000001011000011100000001000000110000111000;  // Label: 5
image_mem[165] = 64'b0011100000110000001110000001110000011000001100000011110000111000;  // Label: 3
image_mem[166] = 64'b0011100001001100010011000011110000000100000001000000110000011000;  // Label: 6
image_mem[167] = 64'b0000110000011000000110000000110000000100000001000000110001111000;  // Label: 5
image_mem[168] = 64'b0000100000001000000110000001100000111100011001000010010000111000;  // Label: 9
image_mem[169] = 64'b0011100000101100001000000010110000110100001001000010110000111000;  // Label: 9
image_mem[170] = 64'b0001100000011100000111000001110000011100001101000011111000011000;  // Label: 8
image_mem[171] = 64'b0001100000011000001111100111011000110100000011000000100000010000;  // Label: 4
image_mem[172] = 64'b0011100000001100000011000000100000011000000101000001110000011000;  // Label: 2
image_mem[173] = 64'b0001100000011000000111000001110000011100000110000001100000011000;  // Label: 1
image_mem[174] = 64'b0011110000100100001000000001110000001000000100000001010000011100;  // Label: 3
image_mem[175] = 64'b0000100000001000000100000001110001111100001000000011100000111000;  // Label: 7
image_mem[176] = 64'b0000100000001000000100000011100000010000001100000011110000011000;  // Label: 7
image_mem[177] = 64'b0000110001111100001110000001100000010000000100000001110000001100;  // Label: 2
image_mem[178] = 64'b0001110000111100000010000001100000010000000100000001010000011100;  // Label: 2
image_mem[179] = 64'b0011110000110000011000000011100000011000000100000011010000011100;  // Label: 3
image_mem[180] = 64'b0001000000101100001000000010000000111100001001000010010000110000;  // Label: 9
image_mem[181] = 64'b0011100000100100001011000001100000110100001001000010010000011000;  // Label: 8
image_mem[182] = 64'b0001110000110100001001000010010000100100001001000010110000011100;  // Label: 0
image_mem[183] = 64'b0001110000110000001100000001000000011000001100000011010000011100;  // Label: 3
image_mem[184] = 64'b0001110000111100000011000000100000011000001100000011110000011000;  // Label: 2
image_mem[185] = 64'b0011100011111000001100000011000000100000001000000011100000011000;  // Label: 2
image_mem[186] = 64'b0001110000110000001100000011000000011100000001000001110000111100;  // Label: 5
image_mem[187] = 64'b0011100001101100010011000011110000000100000001000000100000011000;  // Label: 6
image_mem[188] = 64'b0011110001100100010000000010000000111100001101000011010000011100;  // Label: 9
image_mem[189] = 64'b0001100000100000001000000010000000101100001100100010010000111000;  // Label: 9
image_mem[190] = 64'b0000100000011000000111000011111000100110000001000000110000001000;  // Label: 4
image_mem[191] = 64'b0001100000011000000111000001110000011100000110000001100000011000;  // Label: 1
image_mem[192] = 64'b0001110000011000000111000000011000000010000000100001111000111000;  // Label: 5
image_mem[193] = 64'b0001100000010000001100000011110001111100011011000001100000010000;  // Label: 4
image_mem[194] = 64'b0111110000011100000001000000110000011000000100000001111000011100;  // Label: 2
image_mem[195] = 64'b0011110001100100010000000110000000110000001101000011110000111100;  // Label: 3
image_mem[196] = 64'b0111000001101100010011000010110000111100000011000001100000010000;  // Label: 6
image_mem[197] = 64'b0001100000011000000100000001110000110110011001000000100000010000;  // Label: 4
image_mem[198] = 64'b0001100000111100001101000001110000011100001111000011110000011000;  // Label: 8
image_mem[199] = 64'b0001110000100100001000000010000000011100000001000000010000111100;  // Label: 5
image_mem[200] = 64'b0011110000100000001000000011000000111100001011000010110000011100;  // Label: 9
image_mem[201] = 64'b0001100000110000001000000011010000011110000001100010110000111000;  // Label: 5
image_mem[202] = 64'b0000100000010000000100000011100001110000001000000111110001110000;  // Label: 7
image_mem[203] = 64'b0001100000111100001110000001100000011000001110000010110000001000;  // Label: 8
image_mem[204] = 64'b0011100000111100001000000010100000111100001101000001110000011000;  // Label: 9
image_mem[205] = 64'b0001100000011000000111100111111000110100001001000000100000001000;  // Label: 4
image_mem[206] = 64'b0111100000100100001001000001100000011000001011000010110000011000;  // Label: 8
image_mem[207] = 64'b0011100000011000000110000001100000011000000110000001100000011000;  // Label: 1
image_mem[208] = 64'b0000110000011000001100000011000000011110000001000000110001111100;  // Label: 5
image_mem[209] = 64'b0001000000011100001111100011011000100100001011000100100000010000;  // Label: 4
image_mem[210] = 64'b0001100000010000001111000011110000100100000011000000100000010000;  // Label: 4
image_mem[211] = 64'b0001100000110100001000000010100000111100001101000011110000001000;  // Label: 9
image_mem[212] = 64'b0011100001100100010001000011110000000100000001000000110000001000;  // Label: 6
image_mem[213] = 64'b0001100000001100000011000001110000011000001110000011100000011000;  // Label: 1
image_mem[214] = 64'b0001110000100100001001000001100000111000000101000001010000001100;  // Label: 8
image_mem[215] = 64'b0011100001001100011001000011110000000100000001000000100000011000;  // Label: 6
image_mem[216] = 64'b0001100000111100011011000010010000100100001011000011110000011000;  // Label: 0
image_mem[217] = 64'b0001100000010000000100000011110001111100010011000000100000011000;  // Label: 4
image_mem[218] = 64'b0001110000010000000110000000110000000110000001100001110000111100;  // Label: 5
image_mem[219] = 64'b0011110000111100000011000001100000010000000101100001110000011100;  // Label: 2
image_mem[220] = 64'b0000110000001000000010000011110001111000001000000010110000111100;  // Label: 7
image_mem[221] = 64'b0011000000110000001111000111110000111000000110000001000000110000;  // Label: 4
image_mem[222] = 64'b0011000001101100001001000001110000000100000011000001100000011000;  // Label: 6
image_mem[223] = 64'b0011000000110000001111100010011001100100010010000001100000010000;  // Label: 4
image_mem[224] = 64'b0000011000001100000010000000100000001100000011000011111000111100;  // Label: 5
image_mem[225] = 64'b0011100001101100001111000000110000000100000011000000100000001000;  // Label: 6
image_mem[226] = 64'b0001100000111100001001000010010000101100001011000011110000011000;  // Label: 0
image_mem[227] = 64'b0001110000110000001000000010000000111000001101000011110000111000;  // Label: 3
image_mem[228] = 64'b0111110000001100000010000000100000001000000100000001010000011100;  // Label: 2
image_mem[229] = 64'b0011110000110000001100000001000000011000001100000011000000011100;  // Label: 3
image_mem[230] = 64'b0111100001101100011011000011110000001100000011000001100000011000;  // Label: 6
image_mem[231] = 64'b0000100000001000000011000011100000010000000100000001110000011000;  // Label: 7
image_mem[232] = 64'b0011000000100000001000000010000000100000001111100011100000100000;  // Label: 1
image_mem[233] = 64'b0011100000100100000000000010000000111100000001000000010000011000;  // Label: 5
image_mem[234] = 64'b1111100000111000000100000001100000001000000010000000100000001000;  // Label: 1
image_mem[235] = 64'b0001000000010000000111100111111000010100000110000001100000010000;  // Label: 4
image_mem[236] = 64'b0000110000001000000111000011110000111000000100000001110000011100;  // Label: 7
image_mem[237] = 64'b0011100000101000001001000011110000000100000001000000110000011000;  // Label: 6
image_mem[238] = 64'b0000110000010000000100000000110000001100000101000010010000111100;  // Label: 8
image_mem[239] = 64'b0011100000101100000111000001100000011000001110000011100000011000;  // Label: 8
image_mem[240] = 64'b0001110000100000011000000110000000111110000001000000110000111100;  // Label: 5
image_mem[241] = 64'b0000100000011000000100000000110000001110000001100000110000111000;  // Label: 5
image_mem[242] = 64'b0010000000111100001111000011100000011000000110000001100000011000;  // Label: 1
image_mem[243] = 64'b0001100000110100001001000010010000111100000011000000110000001000;  // Label: 6
image_mem[244] = 64'b0111100000011000000100000001000000110000001001000011110000011000;  // Label: 2
image_mem[245] = 64'b0001100000011100000111000001100000011100001001000010010000111000;  // Label: 8
image_mem[246] = 64'b0001100000100100001001000001110000011100001110000011110000011000;  // Label: 8
image_mem[247] = 64'b0000100000001000000100000011000000111100001001000011110000110000;  // Label: 9
image_mem[248] = 64'b0000110000011000000100000001000000011100001111100011111000111000;  // Label: 9
image_mem[249] = 64'b0000100000011000000100000011110001111000001000000110110000111000;  // Label: 7
image_mem[250] = 64'b0001100000101000010011000100110000111100000010000000100000001000;  // Label: 6
image_mem[251] = 64'b0011110000011100000010000001000000010000000100000001111000001100;  // Label: 2
image_mem[252] = 64'b0001110001111100000010000001100000010000000100000001111000011100;  // Label: 2
image_mem[253] = 64'b1111110001011100000110000001000000010000001111000001110000011100;  // Label: 2
image_mem[254] = 64'b0011100000100110001000000011100000011000001000000001010000011100;  // Label: 3
image_mem[255] = 64'b0000100000011000000111000011011000000100000011000000110000001000;  // Label: 4
    end


    integer i;

    initial begin
        $display("[Testbench] Starting simulation");
        rst = 1;
        #40 rst = 0;



        // === Send images one by one and store results ===
        for (i = 0; i < 256; i = i + 1) begin
            image = image_mem[i];

            // Wait until output is ready
            wait (done == 1);
            #500; // wait a few cycles for stability

            predict_result[i] = predict_idx;

            $display("Image[%0d] â Predict = %0d", i, predict_idx);

            // Reset FSM to allow next image (if needed)
            rst = 1;
            #40 rst = 0;

        end

        $display("[Testbench] All images processed");

        // Optional: dump results
        for (i = 0; i < 256; i = i + 1) begin
            $display("Result[%0d] = %0d", i, predict_result[i]);
        end

        $finish;
    end

endmodule